`timescale 1ns / 1ps
module control_unit(
    input [7:0] instruction
    );


endmodule

`timescale 1ns / 1ps

module microprocessor(
    input [7:0] instruction,
    output [3:0] first_segment,
    output [3:0] second_segment
    );


endmodule
